// hello world
$display("lane_data_0=%h", rt_hdmi_if.lane_data_0);
$display("lane_data_1=%h", rt_hdmi_if.lane_data_1);
$display("lane_data_2=%h", rt_hdmi_if.lane_data_2);
$display("lane_data_3=%h", rt_hdmi_if.lane_data_3);
